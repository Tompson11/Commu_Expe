module transmitor(
	input IsTransmit,
	input has_error,
	input sys_clk,
	input reset,
	output signed [3:0] channel_outI,
	output signed [3:0] channel_outQ
);

wire clk_1, clk_2;
wire [3:0] I,Q;
wire [3:0] I_out,Q_out;
wire m_out;
wire [1:0] conv_out;
wire conv_S;

assign channel_outI = I_out & {4{IsTransmit}};
assign channel_outQ = Q_out & {4{IsTransmit}};

ClkGen Cg(
    .sys_clk	(	sys_clk	),
    .reset		(	reset		),
    .clk_1		(	clk_1		),
    .clk_2		(	clk_2		)
  );
  
 M_sequence_gen M(
	.clk(clk_2),
	.m_out(m_out),
	.reset(reset)
	);

conv_code Conv(
	.clk(clk_2),
	.reset(reset),
	.m_out(m_out),
	.conv_out(conv_out)
	);

P_to_S P2S(
	.clk(clk_1),
	.conv_out(conv_out),
	.reset(reset),
	.conv_S(conv_S)
	);

QAM QAM(
	.clk(clk_1),
	.reset(reset),
	.conv_S(conv_S),
	.I(I),
	.Q(Q)
	);

Channel channel(
	.clk(clk_1),
	.reset(reset),
	.has_error(has_error),
	.I_in(I),
	.Q_in(Q),
	.I_out(I_out),
	.Q_out(Q_out)
	);

endmodule